module pref

[heap]
pub struct Preferences {
pub mut:
	path     string
	is_test  bool
	out_name string
}
